`timescale 1ns/100ps

`include "tartcfg.v"

module tart_block_tb;

   //-------------------------------------------------------------------------
   //
   //  Settings.
   //
   //-------------------------------------------------------------------------
   //  Antenna + accumulator settings:
   parameter AXNUM = `NUM_ANTENNA; // Number of antenna inputs
   parameter NSB   = AXNUM-1;
   parameter ACCUM = `ACCUM_BITS;  // Bit-width of the accumulators
   parameter BLOCK = ACCUM;        // Block samples-counter bits
   parameter MSB   = BLOCK-1;      // Accumulator MSB
   parameter TRATE = `TMUX_RATE;   // Time-multiplexing rate
   parameter TBITS = `TMUX_BITS;   // TMUX bits

   //  Settings for the visibilities data banks:
   parameter BREAD = NREAD << 2;
   parameter XBITS = `BANK_BITS; // Bank-counter bit-width; of the b
   parameter XSB   = XBITS-1;    // MSB of the bank-counter

   //  Internal correlator data-bus settings:
   parameter CBITS = `BANK_BITS + `READ_BITS;
   parameter CSB   = CBITS-1;

   //  External Wishbone-like bus setttings:
   parameter ABITS = `WBADR_BITS;  // Address bit-width
   parameter ASB   = ABITS-1;      // Address MSB
   parameter BBITS = `WBBUS_BITS;  // Bit-width for the SoC WB bus
   parameter BSB   = BBITS-1;      // Bus MSB

   parameter COUNT = 8; // count down from:  (1 << COUNT) - 1;
//    parameter COUNT = 9; // count down from:  (1 << COUNT) - 1;
//    parameter COUNT = 12; // count down from:  (1 << COUNT) - 1;

   //  Read-back settings:
//    parameter NREAD = 24;
   parameter NREAD = 96;
//    parameter NREAD = 120;
//    parameter NREAD = `READ_COUNT >> 2;
//    parameter NREAD = `READ_COUNT;

   //  Additional simulation settings:
   parameter RNG   = `RANDOM_DATA; // Use random antenna data?
   parameter DELAY = `DELAY;       // Simulated combinational delay


   //-------------------------------------------------------------------------
   //
   //  Signals.
   //
   //-------------------------------------------------------------------------
   wire [MSB:0] c_dat, c_val, blocksize, checksum;
   wire [CSB:0] c_adr;
   wire [BSB:0] dat, val, drx;
   reg          clk_x = 1, b_clk = 1, rst = 0;
   reg          cyc = 0, stb = 0, we = 0, bst = 0;
   reg [3:0]    adr;
   reg [BSB:0]  dtx;
   reg          set = 0, get = 0, fin = 0;
   wire         dsp_en, stuck, limp, ack;
   wire         c_cyc, c_stb, c_we, c_bst, c_ack;
   reg [NSB:0]  data [0:255];
   reg [31:0]   viz = 32'h0;
   reg [4:0]    log_bsize = COUNT[4:0];
   wire         sw, switch;

   assign dsp_en = vx_enabled;


   //-------------------------------------------------------------------------
   //  Setup correlator and bus clocks, respectively.
   always #`CLK_X  clk_x <= ~clk_x;
   always #`CLK_B  b_clk <= ~b_clk;
//    always #10 b_clk <= ~b_clk;


   //-------------------------------------------------------------------------
   //  Simulate two visibility calculations.
   integer      num = 0;
   integer      ptr = 0;
   initial begin : SIM_BLOCK
      if (COUNT < 7) begin
`ifdef __USE_FAKE_DSP
         $dumpfile ("fake_tb.vcd");
`else
         $dumpfile ("dsp_tb.vcd");
`endif
         $dumpvars;
      end

      //----------------------------------------------------------------------
      $display("\n%12t: TART DSP settings:", $time);
      $display(  "%12t:  TART I/O bus settings:", $time);
      $display(  "%12t:   SPI data-bus bit-width:  \t\t%3d", $time, BBITS);
      $display(  "%12t:   Number of visibilities banks:    \t%3d", $time, XBITS);
      $display(  "%12t:  TART visibilities read-back settings:", $time);
      $display(  "%12t:   Visibility-data address-width:   \t%3d", $time, ABITS);
      $display(  "%12t:   Data prefetch block-size (words):\t%3d", $time, NREAD);
      $display(  "%12t:   Data prefetch block-size (bytes):\t%3d", $time, BREAD);
      $display(  "%12t:  TART correlator settings:", $time);
      $display(  "%12t:   Accumulator bit-width:   \t\t%3d", $time, ACCUM);
      $display(  "%12t:   Correlator bus data-width:       \t%3d", $time, BLOCK);
      $display(  "%12t:   Correlator bus address-width:    \t%3d", $time, CBITS);

      //----------------------------------------------------------------------
      $display("\n%12t: Generating fake antenna data:", $time);
      if (RNG)
        $display("%12t:  (Data is random values)", $time);
      else
        $display("%12t:  (Data is just increasing counter values)", $time);
      for (ptr = 0; ptr < 256; ptr = ptr+1) begin
         if (RNG) data[ptr] <= $random;
         else     data[ptr] <= ptr;
      end

      //----------------------------------------------------------------------
      #20 $display("\n%12t: Issuing RESET.\n", $time);
      #13 rst <= 1; #40 rst <= 0;

      //----------------------------------------------------------------------
      $display("\n%12t: Setting block-size & beginning correlation (bank 0)", $time);
      #40 set <= 1; num <= 1; dtx <= {1'b1, 2'b00, log_bsize}; ptr <= 4'ha;
      while (!fin) #10;

//       //----------------------------------------------------------------------
//       $display("%12t: Beginning data-acquisition (bank 0):", $time);
//       #40 set <= 1; num <= 1; dtx <= 8'h80; ptr <= 4'h7;
//       while (!fin) #10;

      //----------------------------------------------------------------------
      $display("%12t: Switching banks (bank 1)", $time);
      while (!switching) #10;
      while (switching) #10;

      //----------------------------------------------------------------------
      while (!newblock) #10;
      #10 $display("\n%12t: Reading back visibilities (bank 0)", $time);
      #10 get <= 1; num <= BREAD; ptr <= 4'h8;
      while (!fin) #10;

      //----------------------------------------------------------------------
      while (!switching) #10; while (switching) #10;
      $display("\n%12t: Stopping data-correlation (bank 1)", $time);
      #10 set <= 1; num <= 1; dtx <= 8'h00; ptr <= 4'ha;
      while (!fin) #10;

      //----------------------------------------------------------------------
      while (!newblock) #10;
      #10 $display("\n%12t: Reading back visibilities (bank 1)", $time);
      #10 get <= 1; num <= BREAD; ptr <= 4'h8;
      while (!fin) #10;

      //----------------------------------------------------------------------
//       $display("\n%12t: Reading back counts (bank 1):", $time);
//       #80 get <= 1;
//       while (!fin) #10;

      //----------------------------------------------------------------------
      #80 $display("\n%12t: Simulation finished:", $time);
      $finish;
   end


   //-------------------------------------------------------------------------
   //  Exit if the simulation appears to have stalled.
   //-------------------------------------------------------------------------
   parameter LIMIT = 1000 + (1 << COUNT) * 320;

   initial begin : SIM_FAILED
      $display("%12t: Simulation TIMEOUT limit:\t%12d", $time, LIMIT);
      #LIMIT $display ("\nTIMEOUT!\n");
      $finish;
   end // SIM_FAILED

   always @(posedge b_clk)
     if (newblock)
       $display("%12t: New block available.", $time);


   //-------------------------------------------------------------------------
   //  Read back visibility data, from the correlators' registers.
   //-------------------------------------------------------------------------
   wire       cyc_n = cyc && rxd == 1 && ack;
   integer    rxd = 0;

`ifndef __WB_CLASSIC
   always @(posedge b_clk)
     if (rst) bst <= #DELAY 0;
     else if ((set || get) && num > 2) bst <= #DELAY 1;
     else if (bst && num == 2 && !wat) bst <= #DELAY 0;
`endif

   always @(posedge b_clk)
     if (rst) begin
        {fin, get, set} <= #DELAY 0;
        {cyc, stb, we } <= #DELAY 0;
     end
     else if (set) begin
        $display("%12t: write beginning (num = %1d)", $time, num);
        {fin, get, set} <= #DELAY 0;
        {cyc, stb, we } <= #DELAY 7;
     end
     else if (get) begin
        $display("%12t: read beginning (num = %1d)", $time, num);
        {fin, get, set} <= #DELAY 0;
        {cyc, stb, we } <= #DELAY 6;
     end
     else if (cyc) begin
        if (!stb && ack) $display("%12t: transfer ending", $time);
`ifdef __WB_CLASSIC
        {fin, get, set} <= #DELAY { cyc_n, get, set};
        {cyc, stb, we } <= #DELAY {!cyc_n, !cyc_n, we && !cyc_n};
`else
        {fin, get, set} <= #DELAY { cyc_n, get, set};
        {cyc, stb, we } <= #DELAY {!cyc_n, bst || wat, we && !cyc_n};
`endif
     end
     else begin
        {fin, get, set} <= #DELAY 0;
        {cyc, stb, we } <= #DELAY 0;
     end

   always @(posedge b_clk)
     if (set || get) adr <= #DELAY ptr;

`ifdef __WB_CLASSIC
   always @(posedge b_clk)
     if (cyc && stb && ack) num <= #DELAY num - 1;
`else
   always @(posedge b_clk)
     if (cyc && stb && !wat) num <= #DELAY num - 1;
`endif // __WB_CLASSIC

   always @(posedge b_clk)
     if (get || set) rxd <= num;
     else if (cyc && ack) rxd <= #DELAY rxd - 1;

   //-------------------------------------------------------------------------
   // Display the data, and which correlator and register it is from.
   reg [10:0]   adr_r;
   reg [5:0]    ci;
   reg [4:0]    ri;
   reg [3:0]    rdys = 0, vals = 0;
   wire         rdy = cyc && !we && ack;

//    assign dat = |{rdys, rdy} ? drx : 'bz;
//    assign val = |{vals, set} ? dtx : 'bz;
   wire [2:0]   dst = cyc ? adr : 'bz;
   assign val = cyc && we ? dtx : 'bz;
//    assign dat = rdy || (|rdys) && cyc ? drx : 'bz;
   assign dat = rdy || rdys[0] ? drx : 'bz;

   always @(posedge b_clk) begin
      rdys <= #DELAY {rdys[2:0], rdy};
      vals <= #DELAY {vals[2:0], set};
   end

   reg [1:0] rxc = 0;
   always @(posedge b_clk) begin
      adr_r    <= #DELAY rd_adr;
      {ci, ri} <= #DELAY adr_r;
      if (cyc && stb && !we && ack) begin
         rxc <= #DELAY rxc + 1;
         viz = {dat, viz[31:8]};
         if (rxc == 2'b11)
           $display("%12t: Vis = %08x (d: %8d, c: %02x, r:%02x)", $time, viz, viz, ci, ri);
//            $display("%12t: Vis = %08x (c: %02x, r:%02x)", $time, viz, ci, ri);
      end
   end


   //-------------------------------------------------------------------------
   //  Generate fake DRAM contents.
   //-------------------------------------------------------------------------
   wire [NSB:0] data_w = data[data_index[7:0]];
   integer     data_index = 0;
   reg         ready = 0;
   reg         aq_start = 0, aq_done = 1;
   wire        spi_busy, aq_request;
   wire [2:0]  aq_sample_delay;

   always @(posedge b_clk)
     if (rst)
       {aq_done, aq_start} <= #DELAY 2'b10;
     else if (!aq_start && aq_done && aq_enabled)
       {aq_done, aq_start} <= #DELAY 2'b01;
     else if (!aq_done && aq_start && aq_enabled)
       aq_start <= #DELAY 0;
     else
       aq_done  <= #DELAY aq_done ? aq_done : !aq_enabled;

   always @(posedge b_clk)
     if (rst)
       ready <= #DELAY 0;
     else if (aq_start || aq_request)
       ready <= #DELAY 1;
     else
       ready <= #DELAY 0;

   always @(posedge b_clk)
     if (rst)
       data_index <= #DELAY 0;
     else if (aq_request)
       data_index <= #DELAY data_index + 1;
     else
       data_index <= #DELAY data_index;

   //-------------------------------------------------------------------------
   //  Generate fake antenna data, from the fake DRAM contents.
   wire [NSB:0] antenna;
   reg [3:0]  cnt = 0;
   wire [3:0] next_cnt = wrap_cnt ? 0 : cnt + 1 ;
   wire       wrap_cnt = cnt == TRATE-1;
   integer    rd_adr = 0;

   assign antenna = data[rd_adr[7:0]];

   always @(posedge clk_x)
     if (rst) cnt <= #DELAY 0;
     else     cnt <= #DELAY dsp_en ? next_cnt : cnt;

   always @(posedge clk_x)
     if (rst) rd_adr <= #DELAY 0;
     else     rd_adr <= #DELAY dsp_en && wrap_cnt ? rd_adr + 1 : rd_adr;


   //-------------------------------------------------------------------------
   //     
   //     DATA-ACQUISITION CONTROL AND READ-BACK.
   //     
   //-------------------------------------------------------------------------
   wire [BSB:0] s_dat;
   wire [XSB:0] v_blk;
   wire         s_cyc, s_stb, s_we, s_ack;
   reg          wat = 0;
   wire         overflow, newblock, streamed, accessed, available, switching;
   wire         aq_debug_mode, aq_enabled, vx_enabled, overwrite;

   wire         dsp_cyc, dsp_stb, dsp_we, dsp_bst, dsp_ack;
   wire [XSB:0] dsp_blk;
   wire [7:0]   dsp_dat, dsp_val;

   assign dsp_bst = 1'b0;

// `ifdef __WB_CLASSIC
   always @(posedge b_clk)
     wat <= #DELAY stb && bst && !ack;
// `endif


   //-------------------------------------------------------------------------
   //  Hilbert transform to recover imaginaries.
   //-------------------------------------------------------------------------
   fake_hilbert #( .WIDTH(AXNUM) ) HILB0
     (  .clk(clk_x),
        .rst(rst),
        .en(enable),
        .d(antenna),
        .valid(go),
        .strobe(strobe), // `antenna` data is valid
        .re(re),
        .im(im)
        );


   //-------------------------------------------------------------------------
   //  TART bank-switching unit.
   //-------------------------------------------------------------------------
   tart_bank_switch #( .COUNT(BLOCK) ) SW0
     ( .clk_x(clk_x),
       .clk_i(b_clk),
       .rst_i(rst),
       .ce_i (go),
       .strobe_i(strobe),
       .bcount_i(blocksize),
       .swap_x(swap_x),
       .swap_o(switch)
       );


   //-------------------------------------------------------------------------
   //  A single block of 4 correlators, and implemented using the Xilinx DSP48
   //  primitives.
   //-------------------------------------------------------------------------
   //  The configuration file includes the parameters that determine which
   //  antannae connect to each of the correlators.
`include "../include/tart_pairs.v"
   correlator_block_DSP
     #(  .ACCUM (BLOCK),
         .PAIRS0(PAIRS00_00),
         .PAIRS1(PAIRS00_01),
         .PAIRS2(PAIRS00_02),
         .PAIRS3(PAIRS00_03),
         .DELAY (DELAY)
         ) BLOCK0
       ( .clk_x(clk_x),
         .rst(rst),

         .clk_i(b_clk),
         .cyc_i(cyc),
         .stb_i(stb),
         .we_i (1'b0),
         .bst_i(bst),
         .ack_o(ack),
         .adr_i(adr),
         .dat_i({BLOCK{1'bx}}),
         .dat_o(dat),

         .sw_i(swap_x),
         .en_i(go),
         .re_i(re),
         .im_i(im),

         .bank_o(bankindex)
         );


endmodule // tart_block_tb
