module fifo_sdram_fifo_scheduler(
   input rst,

   input spi_start_aq,

   input write_clk,
   input [7:0] status_cnt,
   output reg aq_write_en = 0,
   output reg aq_read_en = 0,
  
   input bb_clk,

   output reg bb_filled=0,

   input cmd_ready,
   output reg cmd_enable = 0,     
   output reg cmd_wr = 0,
   output reg [SDRAM_ADDRESS_WIDTH-2:0] cmd_address  = 0,
   
   //output reg tx_write_en = 0,
   output reg tx_ready_for_first_read=0,
   input [4:0] tx_status_cnt


   );

   parameter SDRAM_ADDRESS_WIDTH = 22;
   parameter BLOCKSIZE = 8'd32;
   parameter FILL_THRESHOLD = (1 << 9)-BLOCKSIZE;

   reg [SDRAM_ADDRESS_WIDTH-2:0] sdram_wr_ptr = 0;
   reg [SDRAM_ADDRESS_WIDTH-2:0] sdram_rd_ptr = 0;

   reg [1:0] Sync_start = 2'b0;
   wire spi_start_aq_int;
   always @(posedge write_clk) Sync_start[0] <= spi_start_aq;   // notice that we use clkB
   always @(posedge write_clk) Sync_start[1] <= Sync_start[0];   // notice that we use clkB
   assign spi_start_aq_int = Sync_start[1];  // new signal synchronized to (=ready to be used in) clkB domain  
   
   always @(posedge write_clk or posedge rst)
      begin
         if (rst) aq_write_en <= 1'b0;
         else if (spi_start_aq_int) aq_write_en <= 1'b1;
      end

   reg [5:0] rcnt = 6'b0;
   reg read_delay = 1'b0;

   parameter AQ_WAITING       = 3'd0;
   parameter AQ_FIFO_TO_SDRAM = 3'd1;
   parameter TX_WRITING       = 3'd2;
   parameter TX_IDLE          = 3'd3;
   parameter FINISHED         = 3'd4;
   
   reg [2:0] tart_state = AQ_WAITING;
   
//   always @(tart_state)
//      begin
//         case (tart_state)
//            AQ_WAITING:       aq_read_en  <= 1'b0;
//            AQ_FIFO_TO_SDRAM: aq_read_en  <= 1'b1;
//            TX_WRITING:       
//            TX_IDLE:          //tx_write_en <= 1'b0;
//            FINISHED:         //tx_write_en <= 1'b0;
//            default:
//               begin
//                 aq_read_en  <= 1'b0;
//                  tx_write_en <= 1'b0;
//               end
//         endcase
//      end

   always @(posedge bb_clk or posedge rst)
      begin
         if (rst)
            begin
               read_delay <= 1'b0;
               sdram_wr_ptr <= 0;
               sdram_rd_ptr <= 0;
               aq_read_en  <= 1'b0;
               aq_read_en  <= 1'b0;
               tart_state <= AQ_WAITING;
            end
         else
            case (tart_state)
               AQ_WAITING:
                  begin
                     if (sdram_wr_ptr >= FILL_THRESHOLD)
                        begin
                           tart_state <= TX_WRITING;
                           aq_read_en  <= 1'b0;
                        end
                     else if (status_cnt >=  BLOCKSIZE)
                        begin
                           tart_state <= AQ_FIFO_TO_SDRAM;
                           aq_read_en  <= 1'b1;
                        end
                  end
               AQ_FIFO_TO_SDRAM:
                  begin
                     if (read_delay == 1'b1)
                        begin
                           if (rcnt == BLOCKSIZE-1)
                              begin
                                 rcnt <= 6'b0;
                                 aq_read_en  <= 1'b0;
                                 tart_state <= AQ_WAITING;
                              end
                           else  if (cmd_enable) cmd_enable <= 0;
                                 else
                                    begin
                                       if (cmd_ready)
                                          begin
                                             cmd_wr <= 1;
                                             cmd_enable <= 1;
                                             cmd_address <= sdram_wr_ptr;
                                             sdram_wr_ptr <= sdram_wr_ptr + 1'b1;
                                             $display("READING FROM BUFFER  no.%d of %d : %d", rcnt, BLOCKSIZE, sdram_wr_ptr);
                                             rcnt <= rcnt + 1'b1;
                                          end
                                    end
                        end
                     else read_delay <= 1'b1;
                  end
               TX_WRITING:
                     begin
                        bb_filled <= 1;
                        if (tx_status_cnt > 5'd15)
                           begin 
                              $display("WRITING2IDLE: TX BUFFER: bb_rd_ptr: %d", sdram_rd_ptr);
                              tart_state <= TX_IDLE;
                              tx_ready_for_first_read <= 1;
                           end
                        else
                           begin
                              if (cmd_enable) cmd_enable <= 0;
                              else if (cmd_ready)
                                      begin
                                         cmd_wr <= 0;
                                         cmd_enable <= 1;
                                         cmd_address <= sdram_rd_ptr;
                                         sdram_rd_ptr <= sdram_rd_ptr + 1'b1;
                                      end
                          end
                     end
               TX_IDLE:
                  begin
                     if (sdram_rd_ptr < FILL_THRESHOLD)
                        begin 
                           if (tx_status_cnt<5'd5) tart_state <= TX_WRITING;
                        end
                     else tart_state <= FINISHED;
                  end
               FINISHED:
                  begin
                     $display("Finished.");
                  end
            endcase
      end  
endmodule
